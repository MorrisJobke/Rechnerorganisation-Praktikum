-------------------------------------------------------------------------------
-- Title      : microcode_rom
-- Project    : CPU-4
-------------------------------------------------------------------------------
-- File       : microcode_rom.vhd
-- Author     : René Oertel
-- Company    : Chemnitz University of Technology
-- Created    : 2010-09-14
-- Last update: 2010-09-15
-- Platform   : Xilinx Spartan-3E
-------------------------------------------------------------------------------
-- Description: - Memory 64x19 bit for the microcode ROM of the 4-bit CPU
-------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY microcode_rom IS

  PORT (
    address  : IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
    data_out : OUT STD_LOGIC_VECTOR(18 DOWNTO 0));
    
END microcode_rom;

ARCHITECTURE A_behav OF microcode_rom IS

  TYPE rom_type IS ARRAY(0 TO 63) OF STD_LOGIC_VECTOR(18 DOWNTO 0);
  CONSTANT rom : rom_type := (
--  % nnnnnnwmibaaabiimmm %
--  % eeeeeerrorrrabpp112 %
--  % xxxxxx e__lh_______ %
--  % tttttt qre__eeclsss %
--  % ______  eneennnd10  %
--  % mmmmmm  q nn  t     %
--  % cccccc              %
--  % 543210              %                    
    B"0000010000000000001", --00-- % FETCH %
    B"0000100101000000001", --01--
    B"0000000000000010001", --02-- % CCF, SCF %
    B"0000000000001010001", --03-- % ADC, NOT, RRC %
    B"0001010000000010001", --04-- % JPC, JPZ %
    B"0001100000000010001", --05--
    B"0000000000000010001", --06--
    B"0010000000000000001", --07-- % JPC, JPZ (carry, zero gesetzt) %
    B"0010010100100000001", --08--
    B"0010100000000010001", --09--
    B"0010110000000000001", --0A--
    B"0011000100010000001", --0B--
    B"0011010000000010001", --0C--
    B"0000000000000001001", --0D--
    B"0011110000000010001", --0E-- % LD (M) %
    B"0100000000000000001", --0F--
    B"0100010100100000001", --10--
    B"0100100000000010001", --11--
    B"0100110000000000001", --12--
    B"0101000100010000001", --13--  
    B"0101010000000010001", --14--  
    B"0101100000000000010", --15--
    B"0101110100001100010", --16--
    B"0000000000000000010", --17--
    B"0110010000000010001", --18-- % STO (M) %
    B"0110100000000000001", --19--
    B"0110110100100000001", --1A--
    B"0111000000000010001", --1B--
    B"0111010000000000001", --1C--
    B"0111100100010000001", --1D--
    B"0111110000000010001", --1E--
    B"1000001000000000100", --1F-- 
    B"1000011100001000100", --20--
    B"0000001000000000100", --21--
    B"0000000000000010000", --22--
    B"0000000000000010000", --23--
    B"0000000000000010000", --24--
    B"0000000000000010000", --25--
    B"0000000000000010000", --26--
    B"0000000000000010000", --27--
    B"0000000000000010000", --28--
    B"0000000000000010000", --29--
    B"0000000000000010000", --2A--
    B"0000000000000010000", --2B--
    B"0000000000000010000", --2C--
    B"0000000000000010000", --2D--
    B"0000000000000010000", --2E--
    B"0000000000000010000", --2F--
    B"0000000000000010000", --30--
    B"0000000000000010000", --31--
    B"0000000000000010000", --32--
    B"0000000000000010000", --33--
    B"0000000000000010000", --34--
    B"0000000000000010000", --35--
    B"0000000000000010000", --36--
    B"0000000000000010000", --37--
    B"0000000000000010000", --38--
    B"0000000000000010000", --39--
    B"0000000000000010000", --3A--
    B"0000000000000010000", --3B--
    B"0000000000000010000", --3C--
    B"0000000000000010000", --3D--
    B"0000000000000010000", --3E--
    B"1111111111111111111"  --3F-- % dummy   %
  );

BEGIN

  data_out <= rom(CONV_INTEGER(address));

END A_behav;
